
module mems_mics (
	clk_clk,
	mems_that_shit_0_conduit_end_pdm,
	mems_that_shit_0_conduit_end_pdm_clk_out,
	reset_reset_n);	

	input		clk_clk;
	input		mems_that_shit_0_conduit_end_pdm;
	output		mems_that_shit_0_conduit_end_pdm_clk_out;
	input		reset_reset_n;
endmodule

// mems_mics.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module mems_mics (
		input  wire  clk_clk,                                  //                          clk.clk
		input  wire  mems_that_shit_0_conduit_end_pdm,         // mems_that_shit_0_conduit_end.pdm
		output wire  mems_that_shit_0_conduit_end_pdm_clk_out, //                             .pdm_clk_out
		output wire  mems_that_shit_0_conduit_end_dec_clk_out, //                             .dec_clk_out
		input  wire  reset_reset_n                             //                        reset.reset_n
	);

	wire         altpll_0_c0_clk;                                  // altpll_0:c0 -> mems_that_shit_0:pdm_clk
	wire         altpll_0_c1_clk;                                  // altpll_0:c1 -> mems_that_shit_0:dec_clk
	wire         mems_that_shit_0_avalon_master_waitrequest;       // mm_interconnect_0:mems_that_shit_0_avalon_master_waitrequest -> mems_that_shit_0:waitrequest
	wire  [31:0] mems_that_shit_0_avalon_master_address;           // mems_that_shit_0:address -> mm_interconnect_0:mems_that_shit_0_avalon_master_address
	wire   [7:0] mems_that_shit_0_avalon_master_writedata;         // mems_that_shit_0:write_data -> mm_interconnect_0:mems_that_shit_0_avalon_master_writedata
	wire         mems_that_shit_0_avalon_master_write;             // mems_that_shit_0:write -> mm_interconnect_0:mems_that_shit_0_avalon_master_write
	wire         mm_interconnect_0_onchip_memory2_0_s2_chipselect; // mm_interconnect_0:onchip_memory2_0_s2_chipselect -> onchip_memory2_0:chipselect2
	wire   [7:0] mm_interconnect_0_onchip_memory2_0_s2_readdata;   // onchip_memory2_0:readdata2 -> mm_interconnect_0:onchip_memory2_0_s2_readdata
	wire  [11:0] mm_interconnect_0_onchip_memory2_0_s2_address;    // mm_interconnect_0:onchip_memory2_0_s2_address -> onchip_memory2_0:address2
	wire         mm_interconnect_0_onchip_memory2_0_s2_write;      // mm_interconnect_0:onchip_memory2_0_s2_write -> onchip_memory2_0:write2
	wire   [7:0] mm_interconnect_0_onchip_memory2_0_s2_writedata;  // mm_interconnect_0:onchip_memory2_0_s2_writedata -> onchip_memory2_0:writedata2
	wire         mm_interconnect_0_onchip_memory2_0_s2_clken;      // mm_interconnect_0:onchip_memory2_0_s2_clken -> onchip_memory2_0:clken2
	wire  [31:0] master_0_master_readdata;                         // mm_interconnect_1:master_0_master_readdata -> master_0:master_readdata
	wire         master_0_master_waitrequest;                      // mm_interconnect_1:master_0_master_waitrequest -> master_0:master_waitrequest
	wire  [31:0] master_0_master_address;                          // master_0:master_address -> mm_interconnect_1:master_0_master_address
	wire         master_0_master_read;                             // master_0:master_read -> mm_interconnect_1:master_0_master_read
	wire   [3:0] master_0_master_byteenable;                       // master_0:master_byteenable -> mm_interconnect_1:master_0_master_byteenable
	wire         master_0_master_readdatavalid;                    // mm_interconnect_1:master_0_master_readdatavalid -> master_0:master_readdatavalid
	wire         master_0_master_write;                            // master_0:master_write -> mm_interconnect_1:master_0_master_write
	wire  [31:0] master_0_master_writedata;                        // master_0:master_writedata -> mm_interconnect_1:master_0_master_writedata
	wire         mm_interconnect_1_onchip_memory2_0_s1_chipselect; // mm_interconnect_1:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire   [7:0] mm_interconnect_1_onchip_memory2_0_s1_readdata;   // onchip_memory2_0:readdata -> mm_interconnect_1:onchip_memory2_0_s1_readdata
	wire  [11:0] mm_interconnect_1_onchip_memory2_0_s1_address;    // mm_interconnect_1:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire         mm_interconnect_1_onchip_memory2_0_s1_write;      // mm_interconnect_1:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire   [7:0] mm_interconnect_1_onchip_memory2_0_s1_writedata;  // mm_interconnect_1:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_1_onchip_memory2_0_s1_clken;      // mm_interconnect_1:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         rst_controller_reset_out_reset;                   // rst_controller:reset_out -> [altpll_0:reset, mems_that_shit_0:reset, mm_interconnect_0:mems_that_shit_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:master_0_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:onchip_memory2_0_reset1_reset_bridge_in_reset_reset, onchip_memory2_0:reset, onchip_memory2_0:reset2, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;               // rst_controller:reset_req -> [onchip_memory2_0:reset_req, onchip_memory2_0:reset_req2, rst_translator:reset_req_in]

	mems_mics_altpll_0 altpll_0 (
		.clk                (clk_clk),                        //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset), // inclk_interface_reset.reset
		.read               (),                               //             pll_slave.read
		.write              (),                               //                      .write
		.address            (),                               //                      .address
		.readdata           (),                               //                      .readdata
		.writedata          (),                               //                      .writedata
		.c0                 (altpll_0_c0_clk),                //                    c0.clk
		.c1                 (altpll_0_c1_clk),                //                    c1.clk
		.areset             (),                               //        areset_conduit.export
		.scandone           (),                               //           (terminated)
		.scandataout        (),                               //           (terminated)
		.locked             (),                               //           (terminated)
		.phasedone          (),                               //           (terminated)
		.phasecounterselect (4'b0000),                        //           (terminated)
		.phaseupdown        (1'b0),                           //           (terminated)
		.phasestep          (1'b0),                           //           (terminated)
		.scanclk            (1'b0),                           //           (terminated)
		.scanclkena         (1'b0),                           //           (terminated)
		.scandata           (1'b0),                           //           (terminated)
		.configupdate       (1'b0)                            //           (terminated)
	);

	mems_mics_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_clk),                       //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                //    clk_reset.reset
		.master_address       (master_0_master_address),       //       master.address
		.master_readdata      (master_0_master_readdata),      //             .readdata
		.master_read          (master_0_master_read),          //             .read
		.master_write         (master_0_master_write),         //             .write
		.master_writedata     (master_0_master_writedata),     //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                               // master_reset.reset
	);

	MEMS_THAT_SHIT #(
		.IDLE              (4'b0000),
		.TRANSMIT          (4'b0101),
		.WAIT_FOR_TRANSMIT (4'b0001),
		.MEM_SIZE          (25'b0000000000001000000000000)
	) mems_that_shit_0 (
		.reset       (rst_controller_reset_out_reset),             //         reset.reset
		.address     (mems_that_shit_0_avalon_master_address),     // avalon_master.address
		.write_data  (mems_that_shit_0_avalon_master_writedata),   //              .writedata
		.waitrequest (mems_that_shit_0_avalon_master_waitrequest), //              .waitrequest
		.write       (mems_that_shit_0_avalon_master_write),       //              .write
		.clock       (clk_clk),                                    //    clock_sink.clk
		.pdm         (mems_that_shit_0_conduit_end_pdm),           //   conduit_end.pdm
		.pdm_clk_out (mems_that_shit_0_conduit_end_pdm_clk_out),   //              .pdm_clk_out
		.dec_clk_out (mems_that_shit_0_conduit_end_dec_clk_out),   //              .dec_clk_out
		.pdm_clk     (altpll_0_c0_clk),                            //       pdm_clk.clk
		.dec_clk     (altpll_0_c1_clk)                             //       dec_clk.clk
	);

	mems_mics_onchip_memory2_0 onchip_memory2_0 (
		.clk         (clk_clk),                                          //   clk1.clk
		.address     (mm_interconnect_1_onchip_memory2_0_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_onchip_memory2_0_s1_write),      //       .write
		.readdata    (mm_interconnect_1_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_onchip_memory2_0_s1_writedata),  //       .writedata
		.reset       (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),               //       .reset_req
		.address2    (mm_interconnect_0_onchip_memory2_0_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_onchip_memory2_0_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_onchip_memory2_0_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_onchip_memory2_0_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_onchip_memory2_0_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_onchip_memory2_0_s2_writedata),  //       .writedata
		.clk2        (clk_clk),                                          //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),                   // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze      (1'b0)                                              // (terminated)
	);

	mems_mics_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                      (clk_clk),                                          //                                    clk_0_clk.clk
		.mems_that_shit_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                   // mems_that_shit_0_reset_reset_bridge_in_reset.reset
		.mems_that_shit_0_avalon_master_address             (mems_that_shit_0_avalon_master_address),           //               mems_that_shit_0_avalon_master.address
		.mems_that_shit_0_avalon_master_waitrequest         (mems_that_shit_0_avalon_master_waitrequest),       //                                             .waitrequest
		.mems_that_shit_0_avalon_master_write               (mems_that_shit_0_avalon_master_write),             //                                             .write
		.mems_that_shit_0_avalon_master_writedata           (mems_that_shit_0_avalon_master_writedata),         //                                             .writedata
		.onchip_memory2_0_s2_address                        (mm_interconnect_0_onchip_memory2_0_s2_address),    //                          onchip_memory2_0_s2.address
		.onchip_memory2_0_s2_write                          (mm_interconnect_0_onchip_memory2_0_s2_write),      //                                             .write
		.onchip_memory2_0_s2_readdata                       (mm_interconnect_0_onchip_memory2_0_s2_readdata),   //                                             .readdata
		.onchip_memory2_0_s2_writedata                      (mm_interconnect_0_onchip_memory2_0_s2_writedata),  //                                             .writedata
		.onchip_memory2_0_s2_chipselect                     (mm_interconnect_0_onchip_memory2_0_s2_chipselect), //                                             .chipselect
		.onchip_memory2_0_s2_clken                          (mm_interconnect_0_onchip_memory2_0_s2_clken)       //                                             .clken
	);

	mems_mics_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                                       (clk_clk),                                          //                                     clk_0_clk.clk
		.master_0_clk_reset_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                   //      master_0_clk_reset_reset_bridge_in_reset.reset
		.onchip_memory2_0_reset1_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                   // onchip_memory2_0_reset1_reset_bridge_in_reset.reset
		.master_0_master_address                             (master_0_master_address),                          //                               master_0_master.address
		.master_0_master_waitrequest                         (master_0_master_waitrequest),                      //                                              .waitrequest
		.master_0_master_byteenable                          (master_0_master_byteenable),                       //                                              .byteenable
		.master_0_master_read                                (master_0_master_read),                             //                                              .read
		.master_0_master_readdata                            (master_0_master_readdata),                         //                                              .readdata
		.master_0_master_readdatavalid                       (master_0_master_readdatavalid),                    //                                              .readdatavalid
		.master_0_master_write                               (master_0_master_write),                            //                                              .write
		.master_0_master_writedata                           (master_0_master_writedata),                        //                                              .writedata
		.onchip_memory2_0_s1_address                         (mm_interconnect_1_onchip_memory2_0_s1_address),    //                           onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                           (mm_interconnect_1_onchip_memory2_0_s1_write),      //                                              .write
		.onchip_memory2_0_s1_readdata                        (mm_interconnect_1_onchip_memory2_0_s1_readdata),   //                                              .readdata
		.onchip_memory2_0_s1_writedata                       (mm_interconnect_1_onchip_memory2_0_s1_writedata),  //                                              .writedata
		.onchip_memory2_0_s1_chipselect                      (mm_interconnect_1_onchip_memory2_0_s1_chipselect), //                                              .chipselect
		.onchip_memory2_0_s1_clken                           (mm_interconnect_1_onchip_memory2_0_s1_clken)       //                                              .clken
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
